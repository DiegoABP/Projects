`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.04.2021 14:16:36
// Design Name: 
// Module Name: SumaTB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SumaTB;
 reg signed [31:0] A;
 reg signed [31:0] B;
 wire signed [31:0] O;
Suma SU(.A(A),.B(B),.out(O));

initial begin
//0.46   0.79
A=32'b00111110111010111000010100011110;B=32'b00111111010010100011110101110000;
#10;A=32'b00111110111010111000010100011110;B=32'b00111111010010100011110101110000;
#10;A=32'b00111110111010111000010100011110;B=32'b00111110111010111000010100011110;
#10;A=32'b00111110100000000000000000000000;B=32'b00111110100000000000000000000000;
#10;A=32'b00111111010010100011110101110000;B=32'b00111110111010111000010100011110;
#10;A=32'b00111111010010100011110101110000;B=32'b00111111010010100011110101110000;
//0.25 0.5
#10;A=32'b00111110100000000000000000000000;B=32'b00111111000000000000000000000000;
#10;A=32'b00111110100000000000000000000000;B=32'b00111111000000000000000000000000;
#10;A=32'b00111110100000000000000000000000;B=32'b00111110100000000000000000000000;
#10;A=32'b00111110100000000000000000000000;B=32'b00111110100000000000000000000000;
#10;A=32'b00111111000000000000000000000000;B=32'b00111111000000000000000000000000;
#10;A=32'b00111111000000000000000000000000;B=32'b00111111000000000000000000000000;
#10; $finish;
end
endmodule
